// utils.vh
// header files that has global variables and constants to be used in the whole system

// include guards
`ifndef utils_
`define utils_

// Start of include contents

`define ROW_LEN 6			// width of an image
`define COL_LEN 6			// width of an image

reg [11:0] image [35:0];


//= {12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF, 12'h_FFF};

`endif //utils_
